library ieee;
use ieee.std_logic_1164.all;


entity test is
end entity;


architecture tb of test is

    signal end_simulation : boolean := true;

    type vl is ('X', '0', '1', 'Z');
    subtype v0z is vl range '0' to 'Z';
    subtype v01 is vl range '0' to '1';

begin

    process (end_simulation)
    begin
        report "v0z'base: v4l";
        report "v0z'left: " & vl'image(v0z'left); -- '0'
        report "vl'left: " & vl'image(vl'left); -- 'X'
        report "v01'right: " & vl'image(v01'right); -- '1'
        report "vl'right: " & vl'image(vl'right); -- 'Z'
        report "integer'high: " & Integer'image(Integer'high); -- 2147483647
        report "v01'high: " & vl'image(v01'high); -- '1'
        report "integer'low: " & Integer'image(Integer'low); -- -2147483648
        report "v01'low: " & vl'image(v01'low); -- '0'
        -- Position of value in base of type.
        report "v01'pos('Z'): " & Integer'image(v01'pos('Z')); -- 3
        report "vl'pos('Z'): " & Integer'image(vl'pos('Z')); -- 3
        -- Value at position in base of type.
        report "v01'val(1): " & vl'image(v01'val(1)); -- '0'
        report "v1'val(3): " & vl'image(vl'val(3)); -- 'Z'
        -- Value after given value in base of type.
        report "v01'succ('0'): " & vl'image(v01'succ('0')); -- '1'
        report "vl'succ('1'): " & vl'image(vl'succ('1')); -- 'Z'
        -- Value before given value in base of type.
        report "v01'pred('1'): " & vl'image(v01'pred('1')); -- '0'
        report "vl'pred('0'): " & vl'image(vl'pred('0')); -- 'X'
    end process;

    end_simulation <= false after 1 ps;
    assert end_simulation
    report "simulation ended"
    severity failure;

end architecture;
