-- TODO: Write test bench using VUnit.
