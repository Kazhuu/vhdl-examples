context lib_context is
    library ieee;
    use ieee.std_logic_1164.all;
    use test_lib.all;
end context;
