library test_lib;
context test_lib.lib_context;


entity test is
end entity;


architecture tb of test is

    signal test : std_logic := '1';
    signal end_simulation : boolean := true;

begin
    -- TODO: Write rest of this here.

end architecture;


