library ieee;
use ieee.std_logic_1164.all;


entity shift_and_add_multiplier is

end entity;


architecture rtl of shift_and_add_multiplier is

begin

end architecture;
